../modelsim/bubble_sort_moduals/bubble_sort.vhd