../modelsim/bubble_sort_moduals/bubbleSortController.vhd