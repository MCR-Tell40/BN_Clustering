../modelsim/bubble_sort_moduals/sort_function.vhd