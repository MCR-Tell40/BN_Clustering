-- Isolation Flagging count Ram reader